architecture fixed1 of leds is
begin
  (led1, led2, led3, led4, led5) <= std_logic_vector'("00101");
end fixed1;
